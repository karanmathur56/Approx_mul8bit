`timescale 1s / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 29.03.2023 21:52:08
// Design Name: 
// Module Name: approxmul_16bit
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module approxmul_16bit(
    input [7:0] a,b,
    output [15:0] p
    );
    //wire [62:0]w;
    wire [65:1]w;
    
    //D4
//    assign p[0]=a[0]&b[0];
//    assign p[1]=(a[1]&b[0]) | (a[0]&b[1]);
//    assign p[2]=(a[2]&b[0]) | (a[1]&b[1]) | (a[0]&b[2]);
//    assign p[3]=(a[3]&b[0]) | (a[2]&b[1]) | (a[1]&b[2]) | (a[0]&b[3]);
//    assign p[0]=1'b0;
//    assign p[1]=1'b0;
//    assign p[2]=1'b0;
//    assign p[3]=1'b0;
//    assign p[0]=a[0]&b[0];
//    assign p[1]=a[1]&b[0];
//    assign p[2]=a[2]&b[0];
//    assign p[3]=a[3]&b[0];
      assign p[0]=1'b0;
      assign p[1]=1'b1;
      assign p[2]=1'b1;
      assign p[3]=1'b0;
    ha_df ha1((a[4]&b[0]),(a[3]&b[1]),w[1],w[2]);
    ac1 x1((a[5]&b[0]),(a[4]&b[1]),(a[3]&b[2]),(a[2]&b[3]),w[3],w[4]);
    
    ac1 x2((a[6]&b[0]),(a[5]&b[1]),(a[4]&b[2]),(a[3]&b[3]),w[5],w[6]);
    ha_df ha2((a[2]&b[4]),(a[1]&b[5]),w[7],w[8]);
         
    ac2_df y1((a[7]&b[0]),(a[6]&b[1]),(a[5]&b[2]),(a[4]&b[3]),w[9],w[10]);
    ac2_df y2((a[3]&b[4]),(a[2]&b[5]),(a[1]&b[6]),(a[0]&b[7]),w[11],w[12]);
    
    assign w[13] = (a[5]&b[2]) & (a[4]&b[3]);
    assign w[14]=  (a[1]&b[6]) & (a[0]&b[7]);
    
    EC_df z1((a[7]&b[1]),(a[6]&b[2]),(a[5]&b[3]),(a[4]&b[4]),w[13],w[15],w[16],w[17]);
    EC_df z2((a[3]&b[5]),(a[2]&b[6]),(a[1]&b[7]),1'b0,w[14],w[18],w[19],w[20]);
    EC_df z3((a[7]&b[2]),(a[6]&b[3]),(a[5]&b[4]),(a[4]&b[5]),w[15],w[21],w[22],w[23]);
    fa_df fa1((a[3]&b[6]),(a[2]&b[7]),w[18],w[24],w[25]);
    EC_df z4((a[7]&b[3]),(a[6]&b[4]),(a[5]&b[5]),(a[4]&b[6]),w[21],w[26],w[27],w[28]);
    fa_df fa2((a[7]&b[4]),(a[6]&b[5]),w[26],w[29],w[30]);
    
    ac1 x3(w[1],(a[2]&b[2]),(a[1]&b[3]),(a[0]&b[4]),p[4],w[31]); 
    ac1 x4(w[3],w[2],(a[1]&b[4]),(a[0]&b[5]),w[32],w[33]);  
    ac1 x5(w[5],w[7],w[4],(a[0]&b[6]),w[34],w[35]); 
    ac2_df y3(w[9],w[11],w[6],w[8],w[36],w[37]);
    
    //assign w[33]= w[9] | w[11];  //doubt
    assign w[38] = w[9] & w[11]; 
    
    EC_df z5(w[16],w[19],w[10],w[12],w[38],w[39],w[40],w[41]);
    EC_df z6(w[22],w[24],w[17],w[20],w[39],w[42],w[43],w[44]);
    EC_df z7(w[27],w[23],w[25],(a[3]&b[7]),w[42],w[45],w[46],w[47]);
    EC_df z8(w[29],(a[5]&b[6]),(a[4]&b[7]),w[28],w[45],w[48],w[49],w[50]);
    EC_df z9((a[7]&b[5]),(a[6]&b[6]),(a[5]&b[7]),w[30],w[48],w[51],w[52],w[53]);
    fa_df fa3((a[7]&b[6]),(a[6]&b[7]),w[51],w[54],w[55]);
    
    fa_df fa4(w[31],w[32],1'b0,p[5],w[56]);
    fa_df fa5(w[33],w[34],w[56],p[6],w[57]);
    fa_df fa6(w[35],w[36],w[57],p[7],w[58]);
    fa_df fa7(w[37],w[40],w[58],p[8],w[59]);
    fa_df fa8(w[41],w[43],w[59],p[9],w[60]);
    fa_df fa9(w[44],w[46],w[60],p[10],w[61]);
    fa_df fa10(w[49],w[47],w[61],p[11],w[62]);
    fa_df fa11(w[50],w[52],w[62],p[12],w[63]);
    fa_df fa12(w[54],w[53],w[63],p[13],w[64]);
    fa_df fa13((a[7]&b[7]),w[55],w[64],p[14],p[15]);
    //assign p[15]=w[65];

endmodule
